module mips();

control c();

datapath d();

endmodule