module mult3(input [2:0] A, B,
             output [5:0] C);

assign C = A * B;

endmodule