module mult3(a, b, out);

input [2:0] a, b;
output [5:0] c;

assign c = a*b;

endmodule